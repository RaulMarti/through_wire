module through_wire(
    input a,
    output b
);

  assign b = a;
endmodule